// repeat - use to repeat the number of statements for the given number of times.

module repeat_code;
initial begin ;
repeat(4)begin   // Repeat the statements inside 4 times 
  $display ("Good morning");
  $display ("Keep shining");
  $display ("--------------");
end 
end 
endmodule

