teams
c
