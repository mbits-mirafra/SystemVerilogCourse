      10000
      11011
c
