interface adder();
  logic in_a,in_b,in_c;
    logic out_sum,out_carry;
  endinterface
