module AND_Gate(
  input A,
  input B,
  output Y,
  input clk);

  assign Y = A&&B; 
endmodule
