bhavana
Teams
BJT
